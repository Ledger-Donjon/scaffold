-- This file is part of Scaffold
--
-- Scaffold is free software: you can redistribute it and/or modify
-- it under the terms of the GNU Lesser General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.
--
-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU Lesser General Public License for more details.
--
-- You should have received a copy of the GNU Lesser General Public License
-- along with this program.  If not, see <https://www.gnu.org/licenses/>.
--
--
-- Copyright 2025 Ledger SAS, written by Olivier Hériveaux


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.common_pkg.all;


--
-- Configurable ISO14443 module.
--
-- Generates a modulation signal which is fed to an analog front-end (most
-- likely the TRF7970A) and decodes received demodulated sub-carrier signal.
-- Configurable triggers can be generated to synchronize experiments with the RF
-- communication.
--
entity iso14443_module is
port (
    -- System clock.
    clock: in std_logic;
    -- System reset, active low.
    reset_n: in std_logic;
    -- Bus signals
    bus_in: in bus_in_t;

    -- Registers selection signals, from address decoder.
    en_status_control: in std_logic;
    en_config: in std_logic;
    en_data: in std_logic;
    en_timeout: in std_logic;

    -- Output registers
    reg_status: out byte_t;
    reg_data: out byte_t;

    -- 13.56 MHz clock source used for synchronization.
    clock_13_56: in std_logic;
    -- If high, cut RF power (by modulating all the time).
    -- Works for ISO-14443 type A only (requires OOK modulation).
    tearing: in std_logic;

    -- ISO14443 signals
    tx: out std_logic;
    rx: in std_logic;
    trigger: out std_logic );
end;


architecture behavior of iso14443_module is
    -- Status register.
    signal status: byte_t;
    signal busy: std_logic;
    -- Configuration register.
    signal config: byte_t;
    signal trigger_tx_start_en: std_logic;
    signal trigger_tx_end_en: std_logic;
    signal trigger_rx_start_en: std_logic;
    signal trigger_long_en: std_logic;
    signal polarity: std_logic;
    signal use_sync: std_logic;
    -- Timeout register
    signal reg_timeout: std_logic_vector(23 downto 0);

    -- When high, pushes a byte in the FIFO.
    signal push: std_logic;
    -- When high, starts transmitting what has been stored in the FIFO.
    signal start: std_logic;
    -- Triggers generated by the transmit module
    signal trigger_tx_start: std_logic;
    signal trigger_tx_end: std_logic;
    signal trigger_rx_start: std_logic;
    signal trigger_long: std_logic;
    -- Trigger asserted when reception begin.
    signal trigger_rx: std_logic;
    -- High during one clock cycle when a bit has been received.
    signal rx_bit_valid: std_logic;
    -- Received bit value. Valid only if rx_bit_valid is high.
    signal rx_bit_out: std_logic;
    -- Enables RF power, used for tearing.
    signal power_enable: std_logic;

    -- FIFO control signals
    signal rx_fifo_q: std_logic;
    signal rx_fifo_empty: std_logic;
    signal rx_fifo_empty_z: std_logic;
    signal rx_fifo_rdreq: std_logic;
    signal rx_fifo_usedw: std_logic_vector(11 downto 0);
    signal rx_fifo_usedw_z: std_logic_vector(11 downto 0);
    signal trigger_reg: std_logic;
begin
    -- Timeout register
    -- Default value to 2 seconds.
    e_timeout_reg: entity work.module_wide_reg
    generic map (wideness => 3, reset => x"2faf08")
    port map (clock => clock, reset_n => reset_n, en => en_timeout,
        bus_in => bus_in, value => reg_timeout);

    e_iso14443_tx: entity work.iso14443_tx
    port map (
        clock => clock,
        reset_n => reset_n,
        pattern => bus_in.write_data(1 downto 0),
        power_enable => power_enable,
        polarity => polarity,
        push => push,
        start => start,
        busy => busy,
        use_sync => use_sync,
        clock_13_56 => clock_13_56,
        timeout => reg_timeout,
        rx_fifo_q => rx_fifo_q,
        rx_fifo_empty => rx_fifo_empty,
        rx_fifo_rdreq => rx_fifo_rdreq,
        rx_fifo_usedw => rx_fifo_usedw,
        trigger_tx_start => trigger_tx_start,
        trigger_tx_end => trigger_tx_end,
        trigger_rx_start => trigger_rx_start,
        rx => rx,
        tx => tx );

    push <= en_data and bus_in.write;
    start <= en_status_control and bus_in.write and bus_in.write_data(0);

    p_power_enable: process (clock, reset_n)
    begin
        if reset_n = '0' then
            power_enable <= '0';
        elsif rising_edge(clock) then
            if (en_status_control = '1') and (bus_in.write = '1') then
                power_enable <= (power_enable or bus_in.write_data(1)) and (not bus_in.write_data(2));
            else
                power_enable <= power_enable and (not tearing);
            end if;
        end if;
    end process;

    -- Transmission trigger
    p_trigger: process (clock, reset_n)
    begin
        if reset_n = '0' then
            trigger_reg <= '0';
            trigger_long <= '0';
        elsif rising_edge(clock) then
            -- Trigger long is also reset if push is asserted. This is usefull
            -- when no response is received from the card.
            -- We also need to reset the trigger when there is no response: we
            -- AND with busy for that purpose.
            trigger_long <= (trigger_long and busy and (not push)
                    and (not trigger_rx_start))
                or (trigger_tx_start and trigger_tx_start_en)
                or (trigger_tx_end and trigger_tx_end_en);
            trigger_reg <= (trigger_long and trigger_long_en)
                or (trigger_tx_start and trigger_tx_start_en)
                or (trigger_tx_end and trigger_tx_end_en)
                or (trigger_rx_start and trigger_rx_start_en);
        end if;
    end process;

    trigger <= trigger_reg;

    e_config: entity work.module_reg
    generic map (reset => x"00")
    port map (
        clock => clock,
        reset_n => reset_n,
        en => en_config,
        bus_in => bus_in,
        value => config );

    trigger_tx_start_en <= config(0);
    trigger_tx_end_en <= config(1);
    trigger_rx_start_en <= config(2);
    trigger_long_en <= config(3);
    use_sync <= config(6);
    polarity <= config(7);

    status <= "0000000" & busy;
    reg_status <= status;

    rx_fifo_rdreq <= en_data and bus_in.read;

    -- Reading data register pops the FIFO. We want the usedw and empty signals
    -- of the FIFO before the pop operation, so we save them in registers when
    -- data register is read.
    p_fifo_z: process (clock, reset_n) is
    begin
        if reset_n = '0' then
            rx_fifo_usedw_z <= (others => '0');
            rx_fifo_empty_z <= '0';
        elsif rising_edge(clock) then
            if rx_fifo_rdreq then
                rx_fifo_usedw_z <= rx_fifo_usedw;
                rx_fifo_empty_z <= rx_fifo_empty;
            else
                rx_fifo_usedw_z <= rx_fifo_usedw_z;
                rx_fifo_empty_z <= rx_fifo_empty_z;
            end if;
        end if;
    end process;

    reg_data <= rx_fifo_usedw_z(rx_fifo_usedw_z'high
        downto rx_fifo_usedw_z'high - 5) & rx_fifo_empty_z & rx_fifo_q;
end;
